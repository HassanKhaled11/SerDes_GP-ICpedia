package PARAMETERS_pkg ;

parameter CLOCK_PERIOD = 20 ;

endpackage