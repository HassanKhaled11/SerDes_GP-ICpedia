module PMA_RX #(parameter DATA_WIDTH = 10)
				(
					input RX_POS,
					input RX_NEG,
					//input Ser_in,
					input Rst_n,
					input CLK_5G,
					input RxPolarity,
					output [DATA_WIDTH-1:0] Data_out 
					//output K285
				);

////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////
//////////////// 	CDR should be here	   /////////////////
////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////


////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////
//////////////// 	Serial to parallel	   /////////////////
////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////


  Serial_to_Parallel #(.DATA_WIDTH(DATA_WIDTH)) serialToparallel (

      .Recovered_Bit_Clk(CLK_5G),
      .Ser_in(RX_POS),
      .Rst_n(Rst_n),
      .RxPolarity(RxPolarity),
      .Data_Collected(Data_out)  

  );

endmodule 
