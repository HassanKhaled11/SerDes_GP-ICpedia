module assertion_encoding (
    input reg        Bit_Rate_10,
    input reg        Rst,
    input wire       enable_PMA,
    input wire [9:0] data_out,
    input reg        enable,
    input reg  [7:0] data,
    input reg  [3:0] TXDataK
);
  property enable_pma_value;

  endproperty
endmodule
