`timescale 1ns/10ps

package PARAMETERS_pkg ;

parameter CLOCK_PERIOD_10 = 2 ;
parameter CLOCK_PERIOD_TX = 0.2 ;
parameter CLOCK_PERIOD_PCLK = 8 ;
parameter CLOCK_PERIOD_Ref = 10 ;


typedef enum bit {
    negative,
    positive
  } disparity;
endpackage