module CDR
(
   input               d_slicer_in      ,   
   input               p_slicer_in      ,   
   input               d_slicer_n_in    , 
   input               p_slicer_n_in    ,

   output reg [9 : 0]  Code 

); 



endmodule 