interface BFM_if ;


// PORTS


endinterface