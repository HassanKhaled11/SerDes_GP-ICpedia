interface BFM_if ;

// PORTS
 bit   clk ;
 logic [3:0] A;
 logic [3:0] B;
 logic [3:0] out;


endinterface


interface  golden_if;
 bit   clk ;
 logic [3:0] A;
 logic [3:0] B;
 logic [3:0] out;
endinterface 