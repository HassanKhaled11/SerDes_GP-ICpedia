module PMA_RX #(parameter DATA_WIDTH = 10)
				(
					input RX_POS,
					input RX_NEG,
					input Rst_n
					input CLK_5G,
					input RxPolarity,
					output [DATA_WIDTH-1:0] Data_out ,
					//output K285
				);

////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////
//////////////// 	CDR should be here	   /////////////////
////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////


////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////
//////////////// 	Serial to parallel	   /////////////////
////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////

Serial_to_Parallel #(.DATA_WIDTH(DATA_WIDTH)) serialToparallel (
															.Rst_n            (Rst_n),
															.Recovered_Bit_Clk(Recovered_Bit_Clk), // from cdr sampled clk
															.Ser_in           (Ser_in), // from cdr sampled bit
															.RxPolarity       (RxPolarity), // inport
															//.K285             (K285), // out to comma detection
															.Data_to_Decoder  (Data_out) // parallel data to buffer
															);

endmodule 